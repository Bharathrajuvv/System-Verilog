Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Aug 25 07:54 2025
time=0 clk=0 rst=1 d=1 count=x
time=5 clk=1 rst=1 d=1 count=0
time=10 clk=0 rst=0 d=1 count=0
time=15 clk=1 rst=0 d=1 count=1
time=20 clk=0 rst=0 d=1 count=1
time=25 clk=1 rst=0 d=1 count=2
time=30 clk=0 rst=0 d=1 count=2
time=35 clk=1 rst=0 d=1 count=3
time=40 clk=0 rst=0 d=1 count=3
time=45 clk=1 rst=0 d=1 count=4
time=50 clk=0 rst=0 d=1 count=4
time=55 clk=1 rst=0 d=1 count=5
time=60 clk=0 rst=0 d=1 count=5
time=65 clk=1 rst=0 d=1 count=6
time=70 clk=0 rst=0 d=1 count=6
time=75 clk=1 rst=0 d=1 count=7
time=80 clk=0 rst=0 d=1 count=7
time=85 clk=1 rst=0 d=1 count=8
time=90 clk=0 rst=0 d=1 count=8
time=95 clk=1 rst=0 d=1 count=9
time=100 clk=0 rst=0 d=1 count=9
time=105 clk=1 rst=0 d=1 count=10
time=110 clk=0 rst=0 d=0 count=10
time=115 clk=1 rst=0 d=0 count=9
time=120 clk=0 rst=1 d=0 count=9
time=125 clk=1 rst=1 d=0 count=0
time=130 clk=0 rst=0 d=0 count=0
time=135 clk=1 rst=0 d=0 count=15
time=140 clk=0 rst=0 d=0 count=15
time=145 clk=1 rst=0 d=0 count=14
time=150 clk=0 rst=0 d=0 count=14
time=155 clk=1 rst=0 d=0 count=13
time=160 clk=0 rst=0 d=0 count=13
time=165 clk=1 rst=0 d=0 count=12
time=170 clk=0 rst=0 d=0 count=12
time=175 clk=1 rst=0 d=0 count=11
time=180 clk=0 rst=0 d=0 count=11
time=185 clk=1 rst=0 d=0 count=10
time=190 clk=0 rst=0 d=0 count=10
time=195 clk=1 rst=0 d=0 count=9
time=200 clk=0 rst=0 d=0 count=9
time=205 clk=1 rst=0 d=0 count=8
time=210 clk=0 rst=0 d=0 count=8
time=215 clk=1 rst=0 d=0 count=7
time=220 clk=0 rst=0 d=0 count=7
time=225 clk=1 rst=0 d=0 count=6
time=230 clk=0 rst=1 d=0 count=6
time=235 clk=1 rst=1 d=0 count=0
time=240 clk=0 rst=1 d=0 count=0
time=245 clk=1 rst=1 d=0 count=0
$finish called from file "testbench.sv", line 39.
$finish at simulation time                  250
           V C S   S i m u l a t i o n   R e p o r t 
Time: 250 ns
CPU Time:      0.400 seconds;       Data structure size:   0.0Mb
Mon Aug 25 07:54:33 2025
Finding VCD file...
./test.vcd
[2025-08-25 11:54:33 UTC] Opening EPWave...
