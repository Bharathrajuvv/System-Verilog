// Code your testbench here
// or browse Examples
module inc;
  initial begin
    dis();
  end
endmodule

task dis;
  $display("HI BHARATH");
endtask


Output:
Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Oct  3 09:26 2025
HI BHARATH
           V C S   S i m u l a t i o n   R e p o r t 
Time: 0 ns
