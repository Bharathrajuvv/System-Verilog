// Code your design here
module or_gate(output bit [3:0] s);
  initial begin
    s<=4;
  end
endmodule

