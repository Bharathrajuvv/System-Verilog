Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Aug 25 07:52 2025
$time=0,clk=0,rst=1,inf.d=0
$time=5,clk=1,rst=1,inf.d=0
$time=10,clk=0,rst=0,inf.d=1
$time=15,clk=1,rst=0,inf.d=1
$time=20,clk=0,rst=0,inf.d=1
$time=25,clk=1,rst=0,inf.d=1
$time=30,clk=0,rst=0,inf.d=0
$time=35,clk=1,rst=0,inf.d=0
$time=40,clk=0,rst=0,inf.d=1
$time=45,clk=1,rst=0,inf.d=1
$time=50,clk=0,rst=0,inf.d=0
$time=55,clk=1,rst=0,inf.d=0
$time=60,clk=0,rst=0,inf.d=1
$time=65,clk=1,rst=0,inf.d=1
$time=70,clk=0,rst=0,inf.d=1
$time=75,clk=1,rst=0,inf.d=1
$time=80,clk=0,rst=0,inf.d=1
$time=85,clk=1,rst=0,inf.d=1
$time=90,clk=0,rst=0,inf.d=1
$time=95,clk=1,rst=0,inf.d=1
$time=100,clk=0,rst=0,inf.d=1
$time=105,clk=1,rst=0,inf.d=1
$time=110,clk=0,rst=0,inf.d=1
$time=115,clk=1,rst=0,inf.d=1
$finish called from file "testbench.sv", line 30.
$finish at simulation time                  120
           V C S   S i m u l a t i o n   R e p o r t 
Time: 120 ns
CPU Time:      0.360 seconds;       Data structure size:   0.0Mb
Mon Aug 25 07:52:09 2025
Finding VCD file...
./test.vcd
[2025-08-25 11:52:09 UTC] Opening EPW
